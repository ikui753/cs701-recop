--library ieee;
--use ieee.std_logic_1164.all;
--
--use IEEE.numeric_std.all;
--
--use work.recop_types.all;
--use work.various_constants.all;
--
----entity topLevel is 
----port (
----	
----);